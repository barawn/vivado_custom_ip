// convert the 32-bit incoming stream to a 256-bit outgoing stream
// still keep the header, because it's a 16-bit header
// also collapses the tuser[2:1] (CRC/TKEEP) errors
//
// On the output side, expanding to 256 bits means we have 31 tuser
// bits available from the parity bits. 3 of them are used for the
// collapsed start-of-frame, CRC error, and tkeep errors. That leaves
// 28 bits remaining. To keep track of where TLAST occurred, we
// collapse the 32-bit TKEEP into 8 bits: so
//
// tuser[3] = |TKEEP[0 +: 4]
// tuser[4] = |TKEEP[4 +: 4]
// tuser[5] = |TKEEP[8 +: 4]
// tuser[6] = |TKEEP[12 +: 4]
// tuser[7] = |TKEEP[16 +: 4]
// tuser[8] = |TKEEP[20 +: 4]
// tuser[9] = |TKEEP[24 +: 4]
// tuser[10] = |TKEEP[28 +: 4]
//
// tuser[11:30] are still unused.
//
// We don't use interfaces.vh because this gets used in a block diagram
// and the block diagram editor goes nuts with it. WHATEVER.
//
//

module helix_event_frame_32to256(
            input           aclk,
            input           aresetn,
            
            input   [31:0]  s_axis_tdata,
            input           s_axis_tvalid,
            output          s_axis_tready,
            input   [2:0]   s_axis_tuser,
            input           s_axis_tlast,

            output  [255:0] m_axis_tdata,
            output          m_axis_tvalid,
            input           m_axis_tready,
            output  [10:0]  m_axis_tuser,
            output          m_axis_tlast
    );

    // define interface convenience macros
    `define DEFINE_AXI4S_MIN_IF( prefix , width )                   \
        wire [ width - 1:0] prefix``tdata;                          \
        wire prefix``tvalid;                                        \
        wire prefix``tready
    `define CONNECT_AXI4S_MIN_IF( port_prefix , if_prefix )         \
        .``port_prefix``tdata ( if_prefix``tdata ),                 \
        .``port_prefix``tvalid ( if_prefix``tvalid ),               \
        .``port_prefix``tready ( if_prefix``tready )

    // custom width converter tuser input
    wire [3:0] width_converter_tuser = { 1'b0, s_axis_tuser };
    
    // connection from width converter to register slice
    `DEFINE_AXI4S_MIN_IF(width_to_slice_ , 256);
    // we pick up tkeep here, but it gets collapsed into groups of 4 and shoved into spare tuser bits
    wire    [31:0]  width_to_slice_tkeep;
    // tlast
    wire width_to_slice_tlast;
    // full-width tuser output (4*8 = 32 tuser bits)
    wire [31:0] width_to_slice_tuser_full;
    // vectorized full tuser output. This is an array of 3 8-bit vectors
    wire [7:0] width_to_slice_tuser_vect[3:0];
    // vectorize
    generate
        genvar i,j;
        for (i=0;i<4;i=i+1) begin : VECT_OUTER
            for (j=0;j<8;j=j+1) begin : VECT_INNER
                // i.e. for vect[0] this is 0,4,8,12,16,24,28 (in reverse order obviously)
                assign width_to_slice_tuser_vect[i][j] = width_to_slice_tuser_full[4*j+i];
            end
        end
    endgenerate            
    // generate the register slice's tuser, which has 11 tuser bits.
    // The bottom three tuser bits are compressed along the byte axis (if any of the 8 bits goes, this goes)
    // the top tuser bit coming out of the width converter is always zero, so we don't bother with it here, it'll get optimized away anyway
    // the remaining 8 tuser bits are generated by collapsing tkeep, which is always set in groups of 4 anyway. 
    wire [10:0] width_to_slice_tuser = {|width_to_slice_tkeep[28 +: 4],
                                        |width_to_slice_tkeep[24 +: 4],
                                        |width_to_slice_tkeep[20 +: 4],
                                        |width_to_slice_tkeep[16 +: 4],
                                        |width_to_slice_tkeep[12 +: 4],
                                        |width_to_slice_tkeep[8 +: 4],
                                        |width_to_slice_tkeep[4 +: 4],
                                        |width_to_slice_tkeep[0 +: 4],
                                        |width_to_slice_tuser_vect[2],
                                        |width_to_slice_tuser_vect[1],
                                        |width_to_slice_tuser_vect[0] };
    
    helix_event_frame_resizer u_resizer( .aclk(aclk),.aresetn(aresetn),
                                        `CONNECT_AXI4S_MIN_IF( s_axis_ , s_axis_ ),
                                        .s_axis_tuser(width_converter_tuser),
                                        .s_axis_tlast(s_axis_tlast),
                                        `CONNECT_AXI4S_MIN_IF( m_axis_ , width_to_slice_ ),
                                        .m_axis_tkeep( width_to_slice_tkeep),
                                        .m_axis_tuser( width_to_slice_tuser_full ),
                                        .m_axis_tlast( width_to_slice_tlast));

    // register slice to isolate the collapse logic
    axis_data256_tuser11_pipeline u_slice( .aclk(aclk), .aresetn(aresetn),
                                        `CONNECT_AXI4S_MIN_IF( s_axis_ , width_to_slice_ ),
                                        .s_axis_tuser( width_to_slice_tuser ),
                                        .s_axis_tlast( width_to_slice_tlast ),
                                        `CONNECT_AXI4S_MIN_IF( m_axis_ , m_axis_ ),
                                        .m_axis_tuser(m_axis_tuser),
                                        .m_axis_tlast(m_axis_tlast));                                        
    
endmodule

